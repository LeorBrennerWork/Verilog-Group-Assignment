//yinon zadok
`default_nettype none 
`timescale 1 ns / 1 ps
module KeySchedule_top_level(


);